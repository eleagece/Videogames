library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-------------------------------------------------------------------------------------------------------
-- Entity memoria
-------------------------------------------------------------------------------------------------------
entity memoria is
	port ( clk: in std_logic;
			 e: in std_logic; -- escribir 1
			 dataIn: in std_logic_vector(8 downto 0); -- valor RGB para meter
			 dataOut: out std_logic_vector(8 downto 0); -- valor RGB para sacar
			 dataOut2: out std_logic_vector(8 downto 0);
			 dir: in std_logic_vector(9 downto 0); -- selecciona una de las 128 posiciones para leer o escribir
			 dir2: in std_logic_vector(9 downto 0) );
end memoria;

-------------------------------------------------------------------------------------------------------
-- Architecture
-------------------------------------------------------------------------------------------------------
architecture Behavioral of memoria is

--> Types, signals
type tipo is array(0 to 1023) of std_logic_vector(8 downto 0);
signal datos: tipo:=( -- linea 1
                     "000000111","000000111","000000111","000000111", -- 0-3
							"000000111","000000111","000000111","000000111", -- 4-7
							"000000111","000000111","000000111","000000111", -- 8-11
							"000000111","000000111","000000111","000000111", -- 12-15
							"000000111","000000111","000000111","000000111", -- 16-19
							"000000111","000000111","000000111","000000111", -- 20-23
							"000000111","000000111","000000111","000000111", -- 24-27
							"000000111","000000111","000000111","000000111", -- 28-31
							"000000111","000000111","000000111","000000111", -- 32-35
							 -- linea 2
							"000000111","000000111","000000111","000000111", -- 36-39
							"000000111","000000111","000000111","000000111", -- 40-43
							"000000111","000000111","000000111","000000111", -- 44-47
							"000000111","000000111","000000111","000000111", -- 48-51
							"000000111","000000111","000000111","000000000", -- 52-55
							"000000111","000000111","000000111","000000111", -- 56-59
							"000000111","000000111","000000111","000000111", -- 60-63
							"000000111","000000111","000000111","000000111", -- 64-67
							"000000111","000000111","000000111","000000111", -- 68-71
							 -- linea 3
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000000", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							 -- linea 4
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000000", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							 -- linea 5
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000000","000000000", -- 
							"000000000","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							 -- linea 6
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000000","000000000", -- 
							"000000000","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							 -- linea 7
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000000","000000000","000000000", -- 
							"000000000","000000000","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							 -- linea 8
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000000","000000000","000000000", -- 
							"000000000","000000000","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", --       
							 -- linea 9
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000000","000000000","000000000", -- 
							"000000000","000000000","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", --  
							 -- linea 10
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000000","000000000","000000000", -- 
							"000000000","000000000","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							 -- linea 11
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000000","000000000","000000000", -- 
							"000000000","000000000","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", --
							 -- linea 12
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000000","000000000","000000000", -- 
							"000000000","000000000","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", --
							 -- linea 13
							"000000111","111000000","111000000","111000000", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000000","000000000","000000000", -- 
							"000000000","000000000","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"111000000","111000000","111000000","000000111", --
							 -- linea 14
							"000000111","111000000","111000000","111000000", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000000","000000000","000000000", -- 
							"000000000","000000000","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"111000000","111000000","111000000","000000111", --
							 -- linea 15
							"000000111","111000000","111000000","111000000", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000000","000000000","000000000", -- 
							"000000000","000000000","000000111","000000000", -- 
							"000000000","000000000","000000000","000000111", -- 
							"000000111","000000111","000000111","000000111", -- 
							"111000000","111000000","111000000","000000111", --
							 -- linea 16
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000111","000000111","000000111", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000111","000000111","000000111","000000111", -- 
							"000000111","000000000","000000000","000000000", -- 
							"000000000","000000000","000000111","000000000", -- 
							"000000000","000000000","000000000","000000111", -- 
							"000000111","000000111","000000111","000000000", -- 
							"000000000","000000000","000000000","000000000", --  
							 -- linea 17
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000111","000000111","000000111", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000111","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000111","000000000", -- 
							"000000000","000000000","000000000","000000111", -- 
							"000000111","000000111","000000111","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							 -- linea 18
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000111","000000111","000000111", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000111","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000111","000000000", -- 
							"000000000","000000000","000000000","000000111", -- 
							"000000111","000000111","000000111","000000000", -- 
							"000000000","000000000","000000000","000000000", --  
							 -- linea 19
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000111","000000111","000000111", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000111","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000111","000000000", -- 
							"000000000","000000000","000000000","000000111", -- 
							"000000111","000000111","000000111","000000000", -- 
							"000000000","000000000","000000000","000000000", --
							 -- linea 20
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000111","000000111","000000111", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000111","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000111","000000000", -- 
							"000000000","000000000","000000000","000000111", -- 
							"000000111","000000111","000000111","000000000", -- 
							"000000000","000000000","000000000","000000000", --
							 -- linea 21
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000111","000000111","000000111", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000111","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000111","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", --
							 -- linea 22
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000111", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000111","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000111","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", --
							 -- linea 23
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000111","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", --
							 -- linea 24
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000111","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							 -- linea 25
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							 -- linea 26
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							 -- linea 27
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							 -- linea 28 (fin de imagen)
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							-- linea extra
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000", -- 
							"000000000","000000000","000000000","000000000"); -- 
							
--> Begin architecture
begin

-->> Process
-->>> Proceso de reseteo, lectura y escritura en memoria
process(e,clk)
begin
	if (clk'event and clk='1') then
		if (e='1') then
			datos(conv_integer(dir2))<=dataIn;
		else
			dataOut<=datos(conv_integer(dir));
			dataOut2<=datos(conv_integer(dir2));
		end if;
	end if;
end process;

end Behavioral;
