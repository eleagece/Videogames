library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-------------------------------------------------------------------------------------------------------
-- Entity vgacore
-------------------------------------------------------------------------------------------------------
entity vgacore is
	port ( reset: in std_logic; -- reset
		    clock: in std_logic; -- reloj de la FPGA a 100 Mhz
			 clkTecl: in std_logic; -- reloj del teclado
			 bitSerie: in std_logic; -- bit que se recibe en serie del teclado, primero el menos significativo
		    hsyncb: inout std_logic; -- horizontal (line) sync
		    vsyncb: out std_logic;	-- vertical (frame) sync
		    rgb: out std_logic_vector(8 downto 0); -- red, green, blue colores
		    angulo7seg: out std_logic_vector(6 downto 0); -- Para mostrar el �ngulo
			 simbAngulo7seg: out std_logic_vector(6 downto 0); -- Para mostrar �
			 leds: out std_logic_vector(9 downto 0) ); -- Para mostrar la fuerza
end vgacore;

-------------------------------------------------------------------------------------------------------
-- Architecture
-------------------------------------------------------------------------------------------------------
architecture vgacore_arch of vgacore is

-- Components -----------------------------------------------------------------------------------------
-->> memoria
component memoria is
	port ( clk: in std_logic;
			 e: in std_logic; -- escribir 1
			 dataIn: in std_logic_vector(8 downto 0); -- valor RGB para meter
			 dataOut: out std_logic_vector(8 downto 0); -- valor RGB para sacar
			 dataOut2: out std_logic_vector(8 downto 0);			
			 dir: in std_logic_vector(9 downto 0); -- selecciona una de las 1023 posiciones para leer o escribir
			 dir2: in std_logic_vector(9 downto 0) ); 
end component memoria;

-->> conversor 7 segmentos
component conv7seg is
	port ( entrada: in std_logic_vector(3 downto 0);
			 salida: out std_logic_vector(6 downto 0) );
end component conv7seg;

-- Types, constants, signals --------------------------------------------------------------------------
-->> vgacore pantalla
signal hcnt: std_logic_vector(8 downto 0); -- horizontal pixel counter
signal vcnt: std_logic_vector(9 downto 0); -- vertical line counter

-->> vgacore reloj pantalla
signal contadorClk: std_logic_vector(1 downto 0); -- contador para dividir la frecuencia del contador interno
signal clk: std_logic; -- reloj de la pantalla (12,5 Mhz)

-->> vgacore reloj telara�a
signal contadorClkTelarana: std_logic_vector(21 downto 0);
signal clkTelarana: std_logic;

-->> vgacore reloj bruma
signal contadorClkBruma: std_logic_vector(24 downto 0);
signal clkBruma: std_logic;

-->> memoria (fondo)
signal re,wr: std_logic;
signal datosIn: std_logic_vector(8 downto 0);
signal datosOut: std_logic_vector(8 downto 0);
signal datosOut2: std_logic_vector(8 downto 0);
signal direccion: std_logic_vector(9 downto 0);
signal direccion2: std_logic_vector(9 downto 0);
type arrayFilas is array(0 to 27) of std_logic_vector(9 downto 0); 
signal filaMem: arrayFilas; -- array que guarda 0, 36, 36+36, 36+36+36... para sacar la posici�n en memoria de cada fila

-->> roms (spiderman, venom, luna, tumba)
type sprite is array(0 to 1151) of std_logic_vector(8 downto 0);
type arraySprite is array(0 to 47) of std_logic_vector(10 downto 0);
signal filaSprite: arraySprite; -- array que guarda 0, 24, 24+24, 24+24+24... para sacar la posici�n en rom de cada fila
signal spiderman: sprite:=( -- linea 1
                           "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
									"000000000","000000000","000000000","000000000","000000000","000000000","000000111","000000111",
									"000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
									 -- linea 2
                           "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
									"000000000","000000000","000000000","000000000","000000000","000000000","000000111","000000111",
									"000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
									 -- linea 3
                           "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000000",
									"111000000","111000000","111000000","111000000","111000000","111000000","000000000","000000111",
									"000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
									 -- linea 4
                           "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000000",
									"111000000","111000000","111000000","111000000","111000000","111000000","000000000","000000111",
									"000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
									 -- linea 5
                           "000000111","000000111","000000111","000000111","000000111","000000111","000000000","111000000",
									"111000000","111000000","111000000","111000000","111000000","111000000","111000000","000000000",
									"000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
									 -- linea 6
                           "000000111","000000111","000000111","000000111","000000111","000000111","000000000","111000000",
									"111000000","111000000","111000000","111000000","111000000","111000000","111000000","000000000",
									"000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",                           
									 -- linea 7
                           "000000111","000000111","000000111","000000111","000000111","000000111","000000000","111000000",
									"111000000","111000000","000000000","111000000","111000000","111000000","111000000","000000000",
									"000000000","000000111","000000111","000000111","000000111","000000111","000000111","000000111",                           
									 -- linea 8
                           "000000111","000000111","000000111","000000111","000000111","000000111","000000000","111000000",
									"111000000","111000000","000000000","111000000","111000000","111000000","111000000","000000000",
									"000000000","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
									 -- linea 9
                           "000000111","000000111","000000111","000000111","000000111","000000000","111000000","111000000",
									"111000000","000000000","111111111","000000000","000000000","111000000","000000000","111111111",
									"000000000","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
									 -- linea 10
                           "000000111","000000111","000000111","000000111","000000111","000000000","111000000","111000000",
									"111000000","000000000","111111111","000000000","000000000","111000000","000000000","111111111",
									"000000000","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
									 -- linea 11
                           "000000111","000000111","000000111","000000111","000000111","000000000","111000000","111000000",
									"111000000","000000000","111111111","111111111","111111111","000000000","111111111","111111111",
									"000000000","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
									 -- linea 12
                           "000000111","000000111","000000111","000000111","000000111","000000000","111000000","111000000",
									"111000000","000000000","111111111","111111111","111111111","000000000","111111111","111111111",
									"000000000","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
									 -- linea 13
                           "000000111","000000111","000000111","000000111","000000111","000000000","111000000","111000000",
									"111000000","000000000","111111111","111111111","111111111","000000000","111111111","111111111",
									"000000000","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
									 -- linea 14
                           "000000111","000000111","000000111","000000111","000000111","000000000","111000000","111000000",
									"111000000","000000000","111111111","111111111","111111111","000000000","111111111","111111111",
									"000000000","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
									 -- linea 15
                           "000000111","000000111","000000111","000000111","000000111","000000000","000000000","111000000",
									"111000000","111000000","000000000","111111111","111111111","000000000","111111111","000000000",
									"000000000","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
									 -- linea 16
                           "000000111","000000111","000000111","000000111","000000111","000000000","000000000","111000000",
									"111000000","111000000","000000000","111111111","111111111","000000000","111111111","000000000",
									"000000000","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
									 -- linea 17
                           "000000111","000000111","000000111","000000111","000000111","000000111","000000000","111000000",
									"111000000","111000000","111000000","000000000","000000000","111000000","000000000","111000000",
									"000000000","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
									 -- linea 18
                           "000000111","000000111","000000111","000000111","000000111","000000111","000000000","111000000",
									"111000000","111000000","111000000","000000000","000000000","111000000","000000000","111000000",
									"000000000","000000111","000000111","000000111","000000111","000000111","000000111","000000111", 
									 -- linea 19
                           "000000111","000000111","000000111","000000111","000000000","000000000","000000000","111000000",
									"000000000","111000000","111000000","111000000","111000000","111000000","111000000","111000000",
									"000000000","000000000","000000000","000000111","000000111","000000111","000000111","000000111",
									 -- linea 20
                           "000000111","000000111","000000111","000000111","000000000","000000000","000000000","111000000",
									"000000000","111000000","111000000","111000000","111000000","111000000","111000000","111000000",
									"000000000","000000000","000000000","000000111","000000111","000000111","000000111","000000111",
									 -- linea 21
                           "000000111","000000111","000000111","000000000","111000000","000000111","000000111","111000000",
									"111000000","000000000","111000000","111000000","111000000","111000000","111000000","000000000",
									"111000000","000000111","111000000","000000000","000000111","000000111","000000111","000000111",
									 -- linea 22
                           "000000111","000000111","000000111","000000000","111000000","000000111","000000111","111000000",
									"111000000","000000000","111000000","111000000","111000000","111000000","111000000","000000000",
									"111000000","000000111","111000000","000000000","000000111","000000111","000000111","000000111",
									 -- linea 23
                           "000000111","000000111","000000111","000000000","111000000","000000111","000000111","000000111",
									"111000000","111000000","000000000","000000000","000000000","000000000","000000000","111000000",
									"000000111","000000111","111000000","000000000","000000111","000000111","000000111","000000111",
									 -- linea 24
                           "000000111","000000111","000000111","000000000","111000000","000000111","000000111","000000111",
									"111000000","111000000","000000000","000000000","000000000","000000000","000000000","111000000",
									"000000111","000000111","111000000","000000000","000000111","000000111","000000111","000000111",
									 -- linea 25
                           "000000111","000000111","000000000","111000000","111000000","000000111","000000111","000000000",
									"111000000","111000000","111000000","000000000","111000000","111000000","111000000","000000000",
									"000000111","000000111","111000000","111000000","000000000","000000111","000000111","000000111",
									 -- linea 26
                           "000000111","000000111","000000000","111000000","111000000","000000111","000000111","000000000",
									"111000000","111000000","111000000","000000000","111000000","111000000","111000000","000000000",
									"000000111","000000111","111000000","111000000","000000000","000000111","000000111","000000111",
									 -- linea 27
                           "000000111","000000111","000000000","111000000","111000000","000000000","000000000","000000000",
									"111000000","111000000","000000000","000000000","000000000","111000000","111000000","000000000",
									"000000000","000000000","111000000","111000000","000000000","000000111","000000111","000000111",
									 -- linea 28
                           "000000111","000000111","000000000","111000000","111000000","000000000","000000000","000000000",
									"111000000","111000000","000000000","000000000","000000000","111000000","111000000","000000000",
									"000000000","000000000","111000000","111000000","000000000","000000111","000000111","000000111",
									 -- linea 29
                           "000000111","000000111","000000000","111000000","111000000","111000000","000000000","000000000",
									"000000111","111000000","111000000","000000000","111000000","111000000","000000111","000000000",
									"000000000","111000000","111000000","111000000","000000000","000000111","000000111","000000111",
									 -- linea 30
                           "000000111","000000111","000000000","111000000","111000000","111000000","000000000","000000000",
									"000000111","111000000","111000000","000000000","111000000","111000000","000000111","000000000",
									"000000000","111000000","111000000","111000000","000000000","000000111","000000111","000000111",
									 -- linea 31
                           "000000111","000000111","000000000","111000000","111000000","111000000","000000000","000000000",
									"000000111","111000000","111000000","111000000","111000000","111000000","000000111","000000000",
									"000000000","111000000","111000000","111000000","000000000","000000111","000000111","000000111",
									 -- linea 32
                           "000000111","000000111","000000000","111000000","111000000","111000000","000000000","000000000",
									"000000111","111000000","111000000","111000000","111000000","111000000","000000111","000000000",
									"000000000","111000000","111000000","111000000","000000000","000000111","000000111","000000111",
									 -- linea 33
                           "000000111","000000111","000000000","111000000","111000000","111000000","000000000","000000000",
									"000000111","000000111","111000000","111000000","111000000","000000111","000000111","000000000",
									"000000000","111000000","111000000","111000000","000000000","000000111","000000111","000000111",
									 -- linea 34
                           "000000111","000000111","000000000","111000000","111000000","111000000","000000000","000000000",
									"000000111","000000111","111000000","111000000","111000000","000000111","000000111","000000000",
									"000000000","111000000","111000000","111000000","000000000","000000111","000000111","000000111",
									 -- linea 35
                           "000000111","000000111","000000111","000000000","000000000","000000000","000000111","000000000",
									"000000111","000000111","111000000","111000000","111000000","000000111","000000111","000000000",
									"000000111","000000000","000000000","000000000","000000111","000000111","000000111","000000111",
									 -- linea 36
                           "000000111","000000111","000000111","000000000","000000000","000000000","000000111","000000000",
									"000000111","000000111","111000000","111000000","111000000","000000111","000000111","000000000",
									"000000111","000000000","000000000","000000000","000000111","000000111","000000111","000000111",
									 -- linea 37
                           "000000111","000000111","000000111","000000111","000000111","000000111","000000000","000000111",
									"000000111","000000111","111000000","111000000","111000000","000000111","000000111","000000111",
									"000000000","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
									 -- linea 38
                           "000000111","000000111","000000111","000000111","000000111","000000111","000000000","000000111",
									"000000111","000000111","111000000","111000000","111000000","000000111","000000111","000000111",
									"000000000","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
									 -- linea 39
                           "000000111","000000111","000000111","000000111","000000111","000000000","111000000","111000000",
									"000000111","000000111","000000111","000000000","000000111","000000111","000000111","000000111",
									"111000000","000000000","000000111","000000111","000000111","000000111","000000111","000000111",
									 -- linea 40
                           "000000111","000000111","000000111","000000111","000000111","000000000","111000000","111000000",
									"000000111","000000111","000000111","000000000","000000111","000000111","000000111","000000111",
									"111000000","000000000","000000111","000000111","000000111","000000111","000000111","000000111",
									 -- linea 41
                           "000000111","000000111","000000111","000000111","000000000","000000000","111000000","111000000",
									"111000000","000000111","000000000","000000111","000000000","000000111","111000000","111000000",
									"111000000","000000000","000000000","000000111","000000111","000000111","000000111","000000111",
									 -- linea 42
                           "000000111","000000111","000000111","000000111","000000000","000000000","111000000","111000000",
									"111000000","000000111","000000000","000000111","000000000","000000111","111000000","111000000",
									"111000000","000000000","000000000","000000111","000000111","000000111","000000111","000000111",
									 -- linea 43
                           "000000111","000000111","000000000","000000000","111000000","111000000","111000000","111000000",
									"111000000","000000000","000000111","000000111","000000111","000000000","111000000","111000000",
									"111000000","111000000","111000000","000000000","000000000","000000111","000000111","000000111",
									 -- linea 44
                           "000000111","000000111","000000000","000000000","111000000","111000000","111000000","111000000",
									"111000000","000000000","000000111","000000111","000000111","000000000","111000000","111000000",
									"111000000","111000000","111000000","000000000","000000000","000000111","000000111","000000111",
									 -- linea 45
                           "000000111","000000000","111000000","111000000","111000000","111000000","111000000","111000000",
									"111000000","000000000","000000111","000000111","000000111","000000000","111000000","111000000",
									"111000000","111000000","111000000","111000000","111000000","000000000","000000111","000000111",
									 -- linea 46
                           "000000111","000000000","111000000","111000000","111000000","111000000","111000000","111000000",
									"111000000","000000000","000000111","000000111","000000111","000000000","111000000","111000000",
									"111000000","111000000","111000000","111000000","111000000","000000000","000000111","000000111",
									 -- linea 47
                           "000000111","000000000","000000000","000000000","000000000","000000000","000000000","000000000",
									"000000000","000000000","000000111","000000111","000000111","000000000","000000000","000000000",
									"000000000","000000000","000000000","000000000","000000000","000000000","000000111","000000111",
									 -- linea 48
                           "000000111","000000000","000000000","000000000","000000000","000000000","000000000","000000000",
									"000000000","000000000","000000111","000000111","000000111","000000000","000000000","000000000",
									"000000000","000000000","000000000","000000000","000000000","000000000","000000111","000000111");
signal venom: sprite:=( -- linea 1
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","000000111","000000000","000000000","000000000","000000111","000000111","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 2
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","000000111","000000000","000000000","000000000","000000111","000000111","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 3
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
						     "000000111","000000000","000000000","000000000","000000000","000000000","000000000","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 4
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
						     "000000111","000000000","000000000","000000000","000000000","000000000","000000000","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 5
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
						     "000000000","000000000","000000000","000000000","000000000","000000000","000000000","000000000",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 6
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
						     "000000000","000000000","000000000","000000000","000000000","000000000","000000000","000000000",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 7
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000000",
						     "000000000","000000000","000000000","000000000","000000000","000000000","111111111","000000000",
							  "000000000","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 8
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000000",
						     "000000000","000000000","000000000","000000000","000000000","000000000","111111111","000000000",
							  "000000000","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 9
                       "000000111","000000111","000000111","000000111","000000111","000000111","111111111","000000000",
						     "000000000","000000000","000000000","000000000","000000000","000000000","111111111","000000000",
							  "000000000","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 10
                       "000000111","000000111","000000111","000000111","000000111","000000111","111111111","000000000",
						     "000000000","000000000","000000000","000000000","000000000","000000000","111111111","000000000",
							  "000000000","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 11
                       "000000111","000000111","000000111","000000111","000000111","000000111","111111111","000000000",
						     "000000000","000000000","000000000","000000000","000000000","111111111","111111111","000000000",
							  "000000000","000000000","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 12
                       "000000111","000000111","000000111","000000111","000000111","000000111","111111111","000000000",
						     "000000000","000000000","000000000","000000000","000000000","111111111","111111111","000000000",
							  "000000000","000000000","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 13
                       "000000111","000000111","000000111","000000111","000000111","000000111","111111111","111111111",
						     "000000000","000000000","000000000","000000000","111111111","111111111","000000000","000000000",
							  "000000000","000000000","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 14
                       "000000111","000000111","000000111","000000111","000000111","000000111","111111111","111111111",
						     "000000000","000000000","000000000","000000000","111111111","111111111","000000000","000000000",
							  "000000000","000000000","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 15
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000000","111111111",
						     "111111111","000000000","111111111","111111111","111111111","000000000","000000000","111111111",
							  "000000000","000000000","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 16
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000000","111111111",
						     "111111111","000000000","111111111","111111111","111111111","000000000","000000000","111111111",
							  "000000000","000000000","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 17
                       "000000111","000000111","000000111","000000111","000000111","000000111","111111111","000000000",
						     "111111111","000000000","111111111","000000000","000000000","000000000","000000000","111111111",
							  "000000000","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 18
                       "000000111","000000111","000000111","000000111","000000111","000000111","111111111","000000000",
						     "111111111","000000000","111111111","000000000","000000000","000000000","000000000","111111111",
							  "000000000","000000111","000000111","000000111","000000111","000000111","000000111","000000111", 
								-- linea 19
                       "000000111","000000111","000000111","000000111","000000111","000000000","111111111","000000000",
						     "000000000","000000000","000000000","000000000","000000000","111111111","111111111","000000000",
							  "000000000","000000000","000000000","000000000","000000111","000000111","000000111","000000111",
								-- linea 20
                       "000000111","000000111","000000111","000000111","000000111","000000000","111111111","000000000",
						     "000000000","000000000","000000000","000000000","000000000","111111111","111111111","000000000",
							  "000000000","000000000","000000000","000000000","000000111","000000111","000000111","000000111",
								-- linea 21
                       "000000111","000000111","000000111","000000111","000000000","000000000","000000000","111111111",
						     "000000000","000000000","000000000","000000000","111111111","000000000","000000000","000000000",
							  "000000000","000000000","000000000","000000000","000000000","000000111","000000111","000000111",
								-- linea 22
                       "000000111","000000111","000000111","000000111","000000000","000000000","000000000","111111111",
						     "000000000","000000000","000000000","000000000","111111111","000000000","000000000","000000000",
							  "000000000","000000000","000000000","000000000","000000000","000000111","000000111","000000111",
								-- linea 23
                       "000000111","000000111","000000111","000000111","000000000","000000000","000000000","000000000",
						     "000000000","111111111","000000000","111111111","000000000","000000000","000000000","000000000",
							  "111111111","000000000","000000000","000000000","000000000","000000111","000000111","000000111",
								-- linea 24
                       "000000111","000000111","000000111","000000111","000000000","000000000","000000000","000000000",
						     "000000000","111111111","000000000","111111111","000000000","000000000","000000000","000000000",
							  "111111111","000000000","000000000","000000000","000000000","000000111","000000111","000000111",
								-- linea 25
                       "000000111","000000111","000000111","000000111","000000000","000000000","000000000","111111111",
						     "000000000","000000000","000000000","000000000","000000000","000000000","000000000","111111111",
							  "000000000","000000000","000000000","000000000","000000000","000000111","000000111","000000111",
								-- linea 26
                       "000000111","000000111","000000111","000000111","000000000","000000000","000000000","111111111",
						     "000000000","000000000","000000000","000000000","000000000","000000000","000000000","111111111",
							  "000000000","000000000","000000000","000000000","000000000","000000111","000000111","000000111",
								-- linea 27
                       "000000111","000000111","000000000","111111111","000000000","000000000","000000000","000000000",
						     "111111111","111111111","111111111","000000000","111111111","111111111","111111111","000000000",
							  "000000000","000000000","000000000","000000000","111111111","000000000","000000111","000000111",
								-- linea 28
                       "000000111","000000111","000000000","111111111","000000000","000000000","000000000","000000000",
						     "111111111","111111111","111111111","000000000","111111111","111111111","111111111","000000000",
							  "000000000","000000000","000000000","000000000","111111111","000000000","000000111","000000111",
								-- linea 29
                       "000000111","000000111","111111111","000000000","000000000","000000000","000000000","000000000",
						     "000000000","000000000","000000000","111111111","000000000","000000000","000000000","111111111",
							  "111111111","000000000","000000000","000000000","000000000","111111111","000000000","000000111",
								-- linea 30
                       "000000111","000000111","111111111","000000000","000000000","000000000","000000000","000000000",
						     "000000000","000000000","000000000","111111111","000000000","000000000","000000000","111111111",
							  "111111111","000000000","000000000","000000000","000000000","111111111","000000000","000000111",
								-- linea 31
                       "000000111","000000111","000000000","000000000","000000000","000000000","000000000","000000000",
						     "111111111","111111111","000000000","111111111","000000000","111111111","111111111","000000000",
							  "000000000","000000000","000000000","000000000","000000000","000000000","000000000","000000111",
								-- linea 32
                       "000000111","000000111","000000000","000000000","000000000","000000000","000000000","000000000",
						     "111111111","111111111","000000000","111111111","000000000","111111111","111111111","000000000",
							  "000000000","000000000","000000000","000000000","000000000","000000000","000000000","000000111",
								-- linea 33
                       "000000111","000000111","000000000","000000000","000000000","000000000","000000000","000000111",
						     "000000000","000000000","111111111","000000000","111111111","000000000","000000000","111111111",
							  "111111111","000000111","000000000","000000000","000000000","000000000","000000000","000000111",
								-- linea 34
                       "000000111","000000111","000000000","000000000","000000000","000000000","000000000","000000111",
						     "000000000","000000000","111111111","000000000","111111111","000000000","000000000","111111111",
							  "111111111","000000111","000000000","000000000","000000000","000000000","000000000","000000111",
								-- linea 35
                       "000000111","000000111","000000111","000000000","000000000","000000000","000000111","000000111",
						     "111111111","111111111","000000000","000000000","000000000","111111111","111111111","000000000",
							  "000000000","000000111","000000111","000000000","000000000","000000000","000000111","000000111",
								-- linea 36
                       "000000111","000000111","000000111","000000000","000000000","000000000","000000111","000000111",
						     "111111111","111111111","000000000","000000000","000000000","111111111","111111111","000000000",
							  "000000000","000000111","000000111","000000000","000000000","000000000","000000111","000000111",
								-- linea 37
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000000",
						     "000000000","000000000","000000000","000000000","000000000","000000000","000000000","000000000",
							  "000000000","000000000","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 38
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000000",
						     "000000000","000000000","000000000","000000000","000000000","000000000","000000000","000000000",
							  "000000000","000000000","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 39
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000000","000000000",
						     "000000000","000000000","000000000","000000000","000000000","000000000","000000000","000000000",
							  "000000000","000000000","000000000","000000111","000000111","000000111","000000111","000000111",
								-- linea 40
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000000","000000000",
						     "000000000","000000000","000000000","000000000","000000000","000000000","000000000","000000000",
							  "000000000","000000000","000000000","000000111","000000111","000000111","000000111","000000111",
								-- linea 41
                       "000000111","000000111","000000111","000000111","000000111","000000000","000000000","000000000",
						     "000000000","000000000","000000000","000000000","000000111","000000000","000000000","000000000",
							  "000000000","000000000","000000000","000000000","000000111","000000111","000000111","000000111",
								-- linea 42
                       "000000111","000000111","000000111","000000111","000000111","000000000","000000000","000000000",
						     "000000000","000000000","000000000","000000000","000000111","000000000","000000000","000000000",
							  "000000000","000000000","000000000","000000000","000000111","000000111","000000111","000000111",
								-- linea 43
                       "000000111","000000111","000000111","000000000","000000000","000000000","000000000","000000000",
						     "000000000","000000000","000000000","000000111","000000111","000000111","000000000","000000000",
							  "000000000","000000000","000000000","000000000","000000000","000000000","000000111","000000111",
								-- linea 44
                       "000000111","000000111","000000111","000000000","000000000","000000000","000000000","000000000",
						     "000000000","000000000","000000000","000000111","000000111","000000111","000000000","000000000",
							  "000000000","000000000","000000000","000000000","000000000","000000000","000000111","000000111",
								-- linea 45
                       "000000111","000000111","000000000","000000000","000000000","000000000","000000000","000000000",
						     "000000000","000000000","000000000","000000111","000000111","000000111","000000000","000000000",
							  "000000000","000000000","000000000","000000000","000000000","000000000","000000000","000000111",
								-- linea 46
                       "000000111","000000111","000000000","000000000","000000000","000000000","000000000","000000000",
						     "000000000","000000000","000000000","000000111","000000111","000000111","000000000","000000000",
							  "000000000","000000000","000000000","000000000","000000000","000000000","000000000","000000111",
								-- linea 47
                       "000000111","000000111","000000000","000000000","000000000","000000000","000000000","000000000",
						     "000000000","000000000","000000000","000000111","000000111","000000111","000000000","000000000",
							  "000000000","000000000","000000000","000000000","000000000","000000000","000000000","000000111",
								-- linea 48
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","000000111","000000000","000000000","000000000","000000111","000000111","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111");
signal luna: sprite:=(  -- linea 1
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","000000111","000000111","111111111","111111111","000000111","000000111","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 2
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","000000111","000000111","111111111","111111111","000000111","000000111","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 3
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
						     "000000111","000000111","111111111","111111111","111111111","111111111","000000111","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 4
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
						     "000000111","111111111","111111111","111111111","111111111","111111111","111111111","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 5
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","111111111",
						     "111111111","111111111","111111111","111111111","111111111","111111111","111111111","111111111",
							  "111111111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 6
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","111111111",
						     "111111111","111111111","111111111","111111111","111111111","111111111","111111111","111111111",
							  "111111111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 7
                       "000000111","000000111","000000111","000000111","000000111","000000111","111111111","110110110",
						     "110110110","110110110","111111111","111111111","111111111","111111111","111111111","111111111",
							  "111111111","111111111","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 8
                       "000000111","000000111","000000111","000000111","000000111","000000111","111111111","110110110",
						     "110110110","110110110","111111111","111111111","111111111","111111111","111111111","111111111",
							  "111111111","111111111","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 9
                       "000000111","000000111","000000111","000000111","111111111","111111111","111111111","111111111",
						     "111111111","111111111","110110110","110110110","110110110","111111111","111111111","111111111",
							  "111111111","111111111","111111111","111111111","000000111","000000111","000000111","000000111",
								-- linea 10
                       "000000111","000000111","000000111","000000111","111111111","111111111","111111111","111111111",
						     "111111111","110110110","110110110","110110110","110110110","110110110","110110110","111111111",
							  "111111111","111111111","111111111","111111111","000000111","000000111","000000111","000000111",
								-- linea 11
                       "000000111","000000111","000000111","000000111","111111111","111111111","111111111","111111111",
						     "110110110","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							  "111111111","111111111","110110110","110110110","000000111","000000111","000000111","000000111",
								-- linea 12
                       "000000111","000000111","000000111","111111111","111111111","110110110","110110110","111111111",
						     "110110110","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							  "111111111","110110110","110110110","110110110","111111111","000000111","000000111","000000111",
								-- linea 13
                       "000000111","000000111","000000111","111111111","111111111","110110110","110110110","111111111",
						     "110110110","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							  "111111111","110110110","110110110","110110110","111111111","000000111","000000111","000000111",
								-- linea 14
                       "000000111","000000111","000000111","111111111","111111111","110110110","110110110","111111111",
						     "110110110","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							  "111111111","110110110","110110110","110110110","111111111","000000111","000000111","000000111",
								-- linea 15
                       "000000111","000000111","111111111","110110110","110110110","110110110","110110110","111111111",
						     "110110110","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							  "111111111","111111111","110110110","110110110","111111111","111111000","000000111","000000111",
								-- linea 16
                       "000000111","000000111","111111111","110110110","110110110","110110110","110110110","111111111",
						     "110110110","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							  "110110110","111111111","111111111","111111111","111111111","111111000","000000111","000000111",
								-- linea 17
                       "000000111","000000111","111111111","110110110","110110110","110110110","110110110","111111111",
						     "110110110","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							  "110110110","110110110","111111111","111111111","111111111","111111000","000000111","000000111",
								-- linea 18
                       "000000111","111111111","111111111","110110110","110110110","110110110","110110110","111111111",
						     "111111111","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							  "110110110","110110110","110110110","111111111","111111111","111111000","111111000","000000111",
								-- linea 19
                       "000000111","111111111","110110110","110110110","110110110","110110110","110110110","111111111",
						     "110110110","110110110","110110110","110110110","110110110","111111111","111111111","110110110",
							  "110110110","110110110","110110110","111111111","111111111","111111111","111111000","000000111",
								-- linea 20
                       "000000111","111111111","110110110","110110110","110110110","110110110","110110110","111111111",
						     "110110110","110110110","110110110","111111111","111111111","111111111","111111111","110110110",
							  "110110110","110110110","110110110","111111111","111111111","111111111","111111000","000000111",
								-- linea 21
                       "000000111","111111111","110110110","110110110","110110110","110110110","110110110","111111111",
						     "110110110","110110110","110110110","111111111","111111111","111111111","111111111","110110110",
							  "110110110","110110110","110110110","111111111","111111111","111111111","111111000","000000111",
								-- linea 22
                       "111111111","111111111","110110110","111111111","111111111","111111111","110110110","110110110",
						     "110110110","111111111","111111111","111111111","111111111","111111111","111111111","110110110",
							  "110110110","110110110","110110110","111111111","111111111","111111111","111111000","111111000",
								-- linea 23
                       "111111111","110110110","110110110","110110110","110110110","111111111","110110110","110110110",
						     "110110110","111111111","111111111","111111111","111111111","111111111","111111111","110110110",
							  "110110110","110110110","110110110","111111111","111111111","111111111","111111111","111111000",
								-- linea 24
                       "111111111","110110110","110110110","110110110","110110110","111111111","110110110","110110110",
						     "110110110","111111111","111111111","111111111","111111111","111111111","111111111","111111111",
							  "110110110","110110110","111111111","111111111","111111111","111111111","111111111","111111000",
								-- linea 25
                       "111111111","110110110","110110110","110110110","110110110","111111111","111111111","111111111",
						     "111111111","111111111","111111111","111111111","111111111","111111111","111111111","111111111",
							  "110110110","110110110","111111111","111111111","111111111","111111111","111111111","111111000",
								-- linea 26
                       "111111111","110110110","110110110","110110110","110110110","111111111","111111111","110110110",
						     "110110110","111111111","111111111","111111111","111111111","111111111","111111111","111111111",
							  "111111111","111111111","111111111","111111111","111111111","111111111","111111111","111111000",
								-- linea 27
                       "111111111","110110110","110110110","110110110","110110110","111111111","111111111","110110110",
						     "110110110","111111111","111111111","111111111","111111111","111111111","111111111","111111111",
							  "111111111","111111111","111111111","111111111","111111111","111111111","111111000","111111000",
								-- linea 28
                       "000000111","110110110","110110110","110110110","110110110","111111111","111111111","110110110",
						     "110110110","111111111","111111111","111111111","111111111","111111111","111111111","111111111",
							  "111111111","111111111","111111111","111111111","111111111","111111111","111111000","000000111",
								-- linea 29
                       "000000111","110110110","110110110","110110110","110110110","111111111","111111111","111111111",
						     "111111111","110110110","110110110","110110110","111111111","111111111","111111111","111111111",
							  "111111111","111111111","111111111","111111111","111111111","111111111","111111000","000000111",
								-- linea 30
                       "000000111","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
						     "111111111","110110110","110110110","110110110","111111111","111111111","111111111","110110110",
							  "110110110","110110110","110110110","111111111","111111111","111111000","111111000","000000111",
								-- linea 31
                       "000000111","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
						     "111111111","110110110","110110110","110110110","111111111","111111111","111111111","110110110",
							  "110110110","110110110","110110110","111111111","111111111","111111000","111111000","000000111",
								-- linea 32
                       "000000111","000000111","111111111","111111111","111111111","110110110","110110110","110110110",
						     "111111111","110110110","110110110","110110110","111111111","111111111","111111111","111111111",
							  "111111111","111111111","111111111","111111111","111111111","111111000","000000111","000000111",
								-- linea 33
                       "000000111","000000111","111111111","111111111","111111111","110110110","110110110","110110110",
						     "111111111","110110110","110110110","110110110","111111111","111111111","111111111","111111111",
							  "111111111","111111111","111111111","111111111","111111111","111111000","000000111","000000111",
								-- linea 34
                       "000000111","000000111","111111111","111111111","111111111","111111111","111111111","111111111",
						     "111111111","110110110","110110110","110110110","111111111","111111111","111111111","111111111",
							  "111111111","111111111","111111111","111111111","111111000","111111000","000000111","000000111",
								-- linea 35
                       "000000111","000000111","000000111","111111111","111111111","111111111","111111111","110110110",
						     "110110110","111111111","111111111","111111111","111111111","111111111","111111111","111111111",
							  "111111111","111111111","111111111","111111111","111111000","000000111","000000111","000000111",
								-- linea 36
                       "000000111","000000111","000000111","111111111","111111111","111111111","110110110","110110110",
						     "110110110","110110110","111111111","111111111","111111111","111111111","111111111","111111111",
							  "111111111","111111111","111111111","111111000","111111000","000000111","000000111","000000111",
								-- linea 37
                       "000000111","000000111","000000111","111111111","111111111","111111111","110110110","110110110",
						     "110110110","110110110","111111111","111111111","111111111","111111111","111111111","111111111",
							  "111111111","111111111","111111111","111111000","111111000","000000111","000000111","000000111",
								-- linea 38
                       "000000111","000000111","000000111","000000111","111111111","111111111","110110110","110110110",
						     "110110110","110110110","111111111","111111111","111111111","111111111","111111111","111111111",
							  "111111111","111111111","111111111","111111000","000000111","000000111","000000111","000000111",
								-- linea 39
                       "000000111","000000111","000000111","000000111","111111111","111111111","110110110","110110110",
						     "110110110","110110110","111111111","111111111","111111111","111111111","111111111","111111111",
							  "111111111","111111111","111111000","111111000","000000111","000000111","000000111","000000111",
								-- linea 40
                       "000000111","000000111","000000111","000000111","111111111","111111111","111111111","110110110",
						     "110110110","111111111","111111111","111111111","111111111","111111111","111111111","111111111",
							  "111111111","111111000","111111000","111111000","000000111","000000111","000000111","000000111",
								-- linea 41
                       "000000111","000000111","000000111","000000111","000000111","000000111","111111111","111111111",
						     "111111111","111111111","111111111","111111111","111111111","111111111","111111111","111111111",
							  "111111000","111111000","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 42
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","111111111",
						     "111111111","111111111","111111111","111111111","111111111","111111111","111111111","111111111",
							  "111111000","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 43
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","111111111",
						     "111111111","111111111","111111111","111111111","111111111","111111111","111111111","111111111",
							  "111111000","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 44
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","111111111",
						     "111111111","111111111","111111111","111111111","111111111","111111000","111111000","111111000",
							  "111111000","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 45
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
						     "000000111","111111111","111111111","111111111","111111111","111111000","111111000","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 46
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
						     "000000111","000000111","111111111","111111111","111111000","111111000","000000111","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 47
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
						     "000000111","000000111","000000111","111111111","111111000","000000111","000000111","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
								-- linea 48
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
						     "000000111","000000111","000000111","111111111","111111000","000000111","000000111","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111");
signal tumba: sprite:=( -- linea 1
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 2
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 3
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 4
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","000000111","110110110","110110110","110110110","110110110","000000111","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 5
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","000000111","110110110","110110110","110110110","110110110","000000111","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 6
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","110110110","110110110","110110110","110110110","110110110","110110110","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 7
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","110110110","110110110","110110110","110110110","110110110","110110110","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 8
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","110110110","110110110","110110110","110110110","110110110","110110110","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 9
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","110110110","110110110","110110110","110110110","110110110","110110110","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 10
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","110110110","110110110","110110110","110110110","110110110","110110110","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 11
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","110110110","110110110","110110110","110110110","110110110","110110110","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 12
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","110110110","110110110","110110110","110110110","110110110","110110110","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 13
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","110110110","110110110","110110110","110110110","110110110","110110110","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 14
                       "000000111","000000111","000000111","110110110","110110110","110110110","110110110","110110110",
							  "110110110","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							  "110110110","110110110","110110110","110110110","110110110","000000111","000000111","000000111",
							   -- linea 15
                       "000000111","000000111","000000111","110110110","110110110","110110110","110110110","110110110",
							  "110110110","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							  "110110110","110110110","110110110","110110110","110110110","000000111","000000111","000000111",
							   -- linea 16
                       "000000111","000000111","110110110","110110110","111111111","111111111","111111111","111111111",
							  "111111111","110110110","110110110","111111111","111111111","110110110","111111111","111111111",
							  "111111111","111111111","111111111","111111111","110110110","110110110","000000111","000000111",
							   -- linea 17
                       "000000111","000000111","110110110","110110110","111111111","111111111","111111111","111111111",
							  "111111111","111111111","110110110","111111111","111111111","110110110","111111111","111111111",
							  "111111111","111111111","111111111","111111111","110110110","110110110","000000111","000000111",
							   -- linea 18
                       "000000111","000000111","110110110","110110110","111111111","111111111","110110110","110110110",
							  "111111111","111111111","110110110","111111111","111111111","110110110","111111111","111111111",
							  "110110110","110110110","111111111","111111111","110110110","110110110","000000111","000000111",
							   -- linea 19
                       "000000111","000000111","110110110","110110110","111111111","111111111","110110110","110110110",
							  "111111111","111111111","110110110","111111111","111111111","110110110","111111111","111111111",
							  "110110110","110110110","111111111","111111111","110110110","110110110","000000111","000000111",
							   -- linea 20
                       "000000111","000000111","110110110","110110110","111111111","111111111","111111111","111111111",
							  "111111111","110110110","110110110","111111111","111111111","110110110","111111111","111111111",
							  "111111111","111111111","111111111","111111111","110110110","110110110","000000111","000000111",
							   -- linea 21
                       "000000111","000000111","110110110","110110110","111111111","111111111","111111111","111111111",
							  "111111111","110110110","110110110","111111111","111111111","110110110","111111111","111111111",
							  "111111111","111111111","111111111","111111111","110110110","110110110","000000111","000000111",
							   -- linea 22
                       "000000111","000000111","110110110","110110110","111111111","111111111","110110110","110110110",
							  "111111111","111111111","110110110","111111111","111111111","110110110","111111111","111111111",
							  "110110110","110110110","110110110","110110110","110110110","110110110","000000111","000000111",
							   -- linea 23
                       "000000111","000000111","110110110","110110110","111111111","111111111","110110110","110110110",
							  "111111111","111111111","110110110","111111111","111111111","110110110","111111111","111111111",
							  "110110110","110110110","110110110","110110110","110110110","110110110","000000111","000000111",
							   -- linea 24
                       "000000111","000000111","110110110","110110110","111111111","111111111","110110110","110110110",
							  "111111111","111111111","110110110","111111111","111111111","110110110","111111111","111111111",
							  "110110110","110110110","110110110","110110110","110110110","110110110","000000111","000000111",
							   -- linea 25
                       "000000111","000000111","000000111","110110110","110110110","110110110","110110110","110110110",
							  "110110110","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							  "110110110","110110110","110110110","110110110","110110110","000000111","000000111","000000111",
							   -- linea 26
                       "000000111","000000111","000000111","110110110","110110110","110110110","110110110","110110110",
							  "110110110","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							  "110110110","110110110","110110110","110110110","110110110","000000111","000000111","000000111",
							   -- linea 27
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","110110110","110110110","110110110","110110110","110110110","110110110","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 28
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","110110110","110110110","110110110","110110110","110110110","110110110","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 29
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","110110110","110110110","110110110","110110110","110110110","110110110","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 30
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","110110110","110110110","110110110","110110110","110110110","110110110","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 31
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","110110110","110110110","110110110","110110110","110110110","110110110","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 32
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","110110110","110110110","110110110","110110110","110110110","110110110","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 33
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","110110110","110110110","110110110","110110110","110110110","110110110","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 34
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","110110110","110110110","110110110","110110110","110110110","110110110","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 35
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","110110110","110110110","110110110","110110110","110110110","110110110","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 36
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","110110110","110110110","110110110","110110110","110110110","110110110","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 37
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","110110110","110110110","110110110","110110110","110110110","110110110","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 38
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","110110110","110110110","110110110","110110110","110110110","110110110","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 39
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","110110110","110110110","110110110","110110110","110110110","110110110","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 40
                       "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							  "000000111","110110110","110110110","110110110","110110110","110110110","110110110","000000111",
							  "000000111","000000111","000000111","000000111","000000111","000000111","000000111","000000111",
							   -- linea 41
                       "000000111","000000111","000000111","110110110","110110110","110110110","110110110","110110110",
							  "110110110","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							  "110110110","110110110","110110110","110110110","110110110","000000111","000000111","000000111",
							   -- linea 42
                       "000000111","000000111","000000111","110110110","110110110","110110110","110110110","110110110",
							  "110110110","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							  "110110110","110110110","110110110","110110110","110110110","000000111","000000111","000000111",
							   -- linea 43
                       "000000111","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							  "110110110","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							  "110110110","110110110","110110110","110110110","110110110","110110110","110110110","000000111",
							   -- linea 44
                       "000000111","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							  "110110110","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							  "110110110","110110110","110110110","110110110","110110110","110110110","110110110","000000111",
							   -- linea 45
                       "000000111","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							  "110110110","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							  "110110110","110110110","110110110","110110110","110110110","110110110","110110110","000000111",
							   -- linea 46
                       "110110110","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							  "110110110","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							  "110110110","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							   -- linea 47
                       "110110110","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							  "110110110","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							  "110110110","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							   -- linea 48
                       "110110110","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							  "110110110","110110110","110110110","110110110","110110110","110110110","110110110","110110110",
							  "110110110","110110110","110110110","110110110","110110110","110110110","110110110","110110110");

-->> se�ales de posici�n de spiderman, venom y la telara�a
signal SPx,SPy: std_logic_vector(8 downto 0);
signal VEx,VEy: std_logic_vector(8 downto 0);
signal TEx,TEy: std_logic_vector(8 downto 0);
signal Lx,Ly: std_logic_vector(8 downto 0);
signal Bx1,By1,Bx2,By2,Bx3,By3: std_logic_vector(8 downto 0);

-->> se�ales que indican cu�ndo se debe dibujar qu�
signal pintaBorde,pintaBruma,pintaLuna,pintaTumbaSP,pintaTumbaVE,pintaTelarana,pintaSpiderman,pintaVenom,pintaMemoria: std_logic;

-->> se�ales de choque
signal choqueLimites,choqueEdificios,choqueEnemy: std_logic;

-->> conversores 7 segmentos
signal entrada7seg,entrada7seg2: std_logic_vector(3 downto 0);
signal salida7seg,salida7seg2: std_logic_vector(6 downto 0);

-->> m�quina de estados
type TEstado is (SReset,S1a,S2a,S3a,S1b,S2b,S3b); 
signal estado,nestado:TEstado;

-->> tiro parab�lico
signal t: std_logic_vector (9 downto 0);
signal velocidadY: std_logic_vector (4 downto 0);
signal velocidadX: std_logic_vector (3 downto 0);

-->> teclado
signal data: std_logic_vector (10 downto 0); -- 11 bits acumulados del flujo recibido por bitSerie
signal contador: std_logic_vector (3 downto 0); -- contador para identificar 11 ciclos
signal dataOk: std_logic_vector(7 downto 0); -- 8 bits que identifican tecla actual
signal dataAnt: std_logic_vector(7 downto 0); -- 8 bits que identifican tecla anterior
signal tecladoValido: std_logic; -- Se�al para indicar que se puede leer el valor del teclado
signal lanza: std_logic; -- Bot�n para lanzar el pl�tano

-------------------------------------------------------------------------------------------------------
-- Begin architecture
-------------------------------------------------------------------------------------------------------
begin

-- Combinacional --------------------------------------------------------------------------------------
angulo7seg<=salida7seg;
simbAngulo7seg<=salida7seg2;
lanza<='0' when (tecladoValido='1' and dataOk="01001010") else '1'; -- la se�al de lanza se activa cuando se pulsa el espacio

-- Generates ------------------------------------------------------------------------------------------
-->> generate que indica la fila por la que se va pintando el fondo
filaMem(0)<=(others=>'0');
gen1: for i in 1 to 27 generate
	filaMem(i)<=filaMem(i-1)+"100100";
end generate gen1;

-->> generate que indica la fila por la que se van pintando spiderman, venom, luna y tumbas
filaSprite(0)<=(others=>'0');
gen2: for i in 1 to 47 generate
	filaSprite(i)<=filaSprite(i-1)+"11000";
end generate gen2;

-- Component port maps --------------------------------------------------------------------------------
-->> memoria
memoriaComp: memoria port map (clock,wr,datosIn,datosOut,datosOut2,direccion,direccion2);

-->> conversores 7 segmentos
conv7segComp: conv7seg port map (entrada7seg,salida7seg);
conv7segComp2: conv7seg port map (entrada7seg2,salida7seg2);

-- Process --------------------------------------------------------------------------------------------
-->> proceso A: aumenta hcnt con cada ciclo de reloj desde 0 a 380 y lo vuelve a 0.
A: process(clk,reset)
begin
	-- reset asynchronously clears pixel counter
	if reset='1' then
		hcnt <= "000000000";
	-- horiz. pixel counter increments on rising edge of dot clk
	elsif (clk'event and clk='1') then
		-- horiz. pixel counter rolls-over after 381 pixels
		if hcnt<380 then
			hcnt <= hcnt + 1;
		else
			hcnt <= "000000000";
		end if;
	end if;
end process;

-->> proceso B: aumenta vcnt con cada ciclo de hsyncb desde 0 a 527 y lo vuelve a 0.
B: process(hsyncb,reset)
begin
	-- reset asynchronously clears line counter
	if reset='1' then
		vcnt <= "0000000000";
	-- vert. line counter increments after every horiz. line
	elsif (hsyncb'event and hsyncb='1') then
		-- vert. line counter rolls-over after 528 lines
		if vcnt<527 then
			vcnt <= vcnt + 1;
		else
			vcnt <= "0000000000";
		end if;
	end if;
end process;

-->> proceso C
C: process(clk,reset)
begin
	-- reset asynchronously sets horizontal sync to inactive
	if reset='1' then
		hsyncb <= '1';
	-- horizontal sync is recomputed on the rising edge of every dot clk
	elsif (clk'event and clk='1') then
		-- horiz. sync is low in this interval to signal start of a new line
		if (hcnt>=291 and hcnt<337) then
			hsyncb <= '0';
		else
			hsyncb <= '1';
		end if;
	end if;
end process;

-->> proceso D
D: process(hsyncb,reset)
begin
	-- reset asynchronously sets vertical sync to inactive
	if reset='1' then
		vsyncb <= '1';
	-- vertical sync is recomputed at the end of every line of pixels
	elsif (hsyncb'event and hsyncb='1') then
		-- vert. sync is low in this interval to signal start of a new frame
		if (vcnt>=490 and vcnt<492) then
			vsyncb <= '0';
		else
			vsyncb <= '1';
		end if;
	end if;
end process;

-->> proceso que consigue el reloj de 12,5 Mhz al que funciona la pantalla
process (reset,clock,contadorClk)
begin
	if (reset='1') then
		contadorClk<="00";
		clk<='0';
	elsif clock'event and clock='1' then
		if (contadorClk="11") then
			clk<=not clk;
			contadorClk<="00";
		else
			contadorClk<=contadorClk+1;
		end if;
	end if;
end process;

-->> proceso que consigue el reloj de la telara�a
process (reset,clock,contadorClkTelarana)
begin
	if (reset='1') then
		contadorClkTelarana<=(others=>'0');
		clkTelarana<='0';
	elsif clock'event and clock='1' then
		if (contadorClkTelarana=2500000) then
			clkTelarana<=not clkTelarana;
			contadorClkTelarana<=(others=>'0');
		else
			contadorClkTelarana<=contadorClkTelarana+1;
		end if;
	end if;
end process;

-->> proceso que consigue el reloj de la bruma
process (reset,clock,contadorClkBruma)
begin
	if (reset='1') then
		contadorClkBruma<=(others=>'0');
		clkBruma<='0';
	elsif clock'event and clock='1' then
		if (contadorClkBruma=25000000) then
			clkBruma<=not clkBruma;
			contadorClkBruma<=(others=>'0');
		else
			contadorClkBruma<=contadorClkBruma+1;
		end if;
	end if;
end process;

-->> Proceso de cambio de estado
process(clk,reset)
begin
	if reset='1' then 
		estado<=SReset;
	elsif clk'event and clk='1' then
		estado<=nestado;
	end if;
end process;

-->> Proceso de gu�a de cambio de estado y de cambio de jugador
process (estado,choqueEdificios,choqueEnemy,choqueLimites,lanza)
begin
	nestado<=estado;
	wr<='0';
	case estado is
		when SReset=> -- estado de reset
			nestado<=S1a;
	 -- estados de jugador 1 (spiderman)
		when S1a=> -- estado de espera de lanzamiento
			if (lanza='0') then
				nestado<=S2a; -- vamos al estado de lanzamiento
			end if;
		when S2a=> -- estado de lanzamiento
			if (choqueEdificios='1') then
				wr<='1';
				nestado<=S1b;
			elsif (choqueEnemy='1') then
				nestado<=S3a;
			elsif (choqueLimites='1') then
				nestado<=S1b;
			end if;
		when S3a=> -- estado de victoria de spiderman
	-- estados jugador 2 (venom)
		when S1b=> -- estado de espera de lanzamiento para j2
			if (lanza='0') then
				nestado<=S2b; -- vamos al estado de lanzamiento
			end if;
		when S2b=> -- estado de lanzamiento
			if (choqueEdificios='1') then
				wr<='1';
				nestado<=S1a;
			elsif (choqueEnemy='1') then
				nestado<=S3b;
			elsif (choqueLimites='1') then
				nestado<=S1a;
			end if;
		when S3b=> -- estado de victoria de venom
		when others=> null;
	end case;			
end process;

-->> Proceso que indica cu�ndo se debe dibujar qu�
process(vcnt,hcnt,estado,TEx,TEy,SPx,SPy,VEx,VEy,Bx1,By1)
begin
	pintaBorde<='0';
	pintaTelarana<='0';
	pintaLuna<='0';
	pintaTumbaSP<='0';
	pintaTumbaVE<='0';
	pintaSpiderman<='0';
	pintaVenom<='0';
	pintaMemoria<='0';
	pintaBruma<='0';
	-- activa pintaBorde (m�s prioritario)
	if ((vcnt=0) and (hcnt>0 and hcnt<289)) xor -- horizontal (1 a 288) en vcnt=0
		((vcnt=449) and (hcnt>0 and hcnt<289)) xor -- horizontal (1 a 288) en vcnt=449
		((vcnt>=0 and vcnt<450) and (hcnt=0)) xor -- vertical (0 a 449) en hcnt=0
		((vcnt>=0 and vcnt<450) and (hcnt=289)) then -- vertical (0 a 449) en hcnt=289
		pintaBorde<='1';
	-- activa pintaTelarana
	elsif (hcnt>=TEx and hcnt<=TEx+7 and vcnt>=TEy and vcnt<=TEy+7 and (estado=S2a or estado=S2b)) then
		pintaTelarana<='1';
	-- activa pintaBruma
	elsif (hcnt>=Bx1 and hcnt<=Bx1+50 and vcnt>=By1 AND vcnt<=By1+3) xor
			(hcnt>=Bx2 and hcnt<=Bx2+100 and vcnt>=By2 AND vcnt<=By2+3) xor
			(hcnt>=Bx3 and hcnt<=Bx3+75 and vcnt>=By3 AND vcnt<=By3+3) then
		pintaBruma<='1';
	-- activa pintaLuna
	elsif (hcnt>=Lx and hcnt<=Lx+23 and vcnt>=Ly and vcnt<=Ly+47) then -- Lx-Lx+23(x) (24px)
		pintaLuna<='1';																 -- Ly-Ly+47(y) (48px)
	-- activa pintaTumbaSP
	elsif (hcnt>=SPx and hcnt<=SPx+23 and vcnt>=SPy and vcnt<=SPy+47 and estado=S3b) then -- SPx-SPx+23(x) (24px)
		pintaTumbaSP<='1';																					  -- SPy-SPy+47(y) (48px)
	-- activa pintaTumbaVE
	elsif (hcnt>=VEx and hcnt<=VEx+23 and vcnt>=VEy and vcnt<=VEy+47 and estado=S3a) then -- VEx-VEx+23(x) (24px)
		pintaTumbaVE<='1';																					  -- VEy-VEy+47(y) (48px)
	-- activa pintaSpiderman
	elsif (hcnt>=SPx and hcnt<=SPx+23 and vcnt>=SPy and vcnt<=SPy+47 and estado/=S3b) then -- SPx-SPx+23(x) (24px)
		pintaSpiderman<='1';													  									-- SPy-SPy+47(y) (48px)
	-- activa pintaVenom
	elsif (hcnt>=VEx and hcnt<=VEx+23 and vcnt>=VEy and vcnt<=VEy+47 and estado/=S3a) then -- VEx-VEx+23(x) (24px)
		pintaVenom<='1';																							-- VEy-VEy+47(y) (48px)
	-- activa pintaMemoria (menos prioritario)
	elsif (vcnt>0 and vcnt<449 and hcnt>0 and hcnt<289) then -- 1-288(x) (288px)
		pintaMemoria<='1';												-- 1-448(y) (448px)
	end if;
end process;

-->> Proceso de dibujado en pantalla de borde, telara�a, spiderman, venom, tumbas, luna y memoria
process (pintaBorde,pintaLuna,pintaTumbaSP,pintaTumbaVE,pintaTelarana,pintaSpiderman,pintaVenom,pintaMemoria,datosOut)
begin	
	direccion<=(others=>'1');
	if (pintaBorde='1') then
		rgb<=(others=>'1');
	elsif (pintaBruma='1') then
		rgb<=(others=>'1');
	elsif (pintaLuna='1') then -- x=32 a x=55, y=32 a y=55
		rgb<=luna(conv_integer( filaSprite(conv_integer(vcnt-Ly)) + (hcnt-Lx) ));
	elsif (pintaTumbaSP='1') then -- x=9 a x=32, y=193 a y=240
		rgb<=tumba(conv_integer( filaSprite(conv_integer(vcnt-SPy)) + (hcnt-SPx) ));
	elsif (pintaTumbaVE='1') then -- x=257 a x=280, y=193 a y=240
		rgb<=tumba(conv_integer( filaSprite(conv_integer(vcnt-VEy)) + (hcnt-VEx) ));
	elsif (pintaSpiderman='1') then -- x=9 a x=32, y=193 a y=240
		rgb<=spiderman(conv_integer( filaSprite(conv_integer(vcnt-SPy)) + (hcnt-SPx) ));
	elsif (pintaVenom='1') then -- x=257 a x=280, y=193 a y=240
		rgb<=venom(conv_integer( filaSprite(conv_integer(vcnt-VEy)) + (hcnt-VEx) ));
	elsif (pintaTelarana='1') then
		rgb<=(others=>'1');
	elsif (pintaMemoria='1') then
		direccion<=filaMem(conv_integer(vcnt(8 downto 4)))+(hcnt(8 downto 3));
		if (datosOut="111000000") then
			rgb<="000000111"; -- el area de impacto se pinta del color de fondo
		else
			rgb<=datosOut; -- pinta en el cuadrado n, la direcci�n de memoria n	
		end if;
	else	
		rgb<=(others=>'0'); 
	end if;
end process;

-->> Proceso de c�lculo de choques
process(datosOut2,TEx,TEy)
begin
	datosIn<="000000111";
	choqueEdificios<='0';
	choqueEnemy<='0';
	choqueLimites<='0';
	direccion2<=filaMem(conv_integer(TEy(8 downto 4)))+(TEx(8 downto 3));
	if (TEx<=0 or TEx>=289 or TEy<=0 or TEy>=449) then
		choqueLimites<='1';
	elsif (datosOut2="000000000" or datosOut2="111111000") then
		choqueEdificios<='1';
	elsif (datosOut2="111000000") then
		choqueEnemy<='1';
	end if;
end process;

-->> Proceso de c�lculo de posici�n de spiderman (y su tumba), venom (y su tumba), luna y telara�a
process(estado,clkTelarana,clkBruma)
begin
	SPx<="000001001"; -- 9 posici�n x desde donde se dibuja a spiderman
	SPy<="011000001"; -- 193 posici�n y desde donde se dibuja a spiderman
	VEx<="100000001"; -- 257 posici�n x desde donde se dibuja a venom
	VEy<="011000001"; -- 193 posici�n y desde donde se dibuja a venom
	Lx<="000100000"; -- 32 posici�n x desde donde se dibuja la luna
	Ly<="000100000"; -- 32 posici�n y desde donde se dibuja la luna
	By1<="000101010";
	By2<="000111111";
	By3<="001100010";
	if (clkBruma'event and clkBruma='1') then
		if (estado=SReset) then
			Bx1<="000000000";
			Bx2<="000001111";
			Bx3<="000010100";
		else
			Bx1<=Bx1+1;
			Bx2<=Bx2+2;
			Bx3<=Bx3+3;
		end if;
	end if;
	if (clkTelarana'event and clkTelarana='1') then
		if ((estado=S1a or estado=S1b) and tecladoValido='1') then 
			-- �ngulo
			if (dataOK="00111000") then -- Pulsa �
				velocidadY<="00000";
				entrada7seg<="0000";
			elsif (dataOK="00110100") then -- Pulsa 1 
				velocidadY<="00001";
				entrada7seg<="0001";
			elsif (dataOK="00111100") then -- Pulsa 2
				velocidadY<="00010";
				entrada7seg<="0010";
			elsif (dataOK="00110010") then -- Pulsa 3
				velocidadY<="00100";
				entrada7seg<="0011";
			elsif (dataOK="01010010") then -- Pulsa 4
				velocidadY<="01000";
				entrada7seg<="0100";
			elsif (dataOK="00111010") then -- Pulsa 5
				velocidadY<="01011";
				entrada7seg<="0101";
			elsif (dataOK="00110110") then -- Pulsa 6
				velocidadY<="01111";
				entrada7seg<="0110";
			elsif (dataOK="01011110") then -- Pulsa 7
				velocidadY<="10000";
				entrada7seg<="0111";
			elsif (dataOK="00111110") then -- Pulsa 8
				velocidadY<="11101";
				entrada7seg<="1000";
			elsif (dataOK="00110001") then -- Pulsa 9
				velocidadY<="10000";
				entrada7seg<="1001";
			elsif (dataOK="01010001") then -- Pulsa 0
				velocidadY<="11100";
				entrada7seg<="1010";
			-- Velocidad
			elsif (dataOK="01001011") then -- Pulsa 1 
				velocidadX<="0001";
				leds<="0000000001";
			elsif (dataOK="00100111") then -- Pulsa 2 
				velocidadX<="0011";
				leds<="0000000011";
			elsif (dataOK="00101111") then -- Pulsa 3
				velocidadX<="0100";
				leds<="0000000111";
			elsif (dataOK="01101011") then -- Pulsa 4
				velocidadX<="0101";
				leds<="0000001111";
			elsif (dataOK="01100111") then -- Pulsa 5
				velocidadX<="0110";
				leds<="0000011111";
			elsif (dataOK="00010111") then -- Pulsa 6
				velocidadX<="0111";
				leds<="0000111111";
			elsif (dataOK="00011011") then -- Pulsa 7
				velocidadX<="1000";
				leds<="0001111111";
			elsif (dataOK="01010111") then -- Pulsa 8
				velocidadX<="1001";
				leds<="0011111111";
			elsif (dataOK="01011111") then -- Pulsa 9
				velocidadX<="1010";
				leds<="0111111111";
			elsif (dataOK="00000111") then -- Pulsa 0
				velocidadX<="1100";
				leds<="1111111111";
			end if;
		end if;
		entrada7seg2<="1111"; -- Para que saque el s�mbolo � (ya no saca una F)
		if (estado=S1a) then
			TEx<=SPx+24;
			TEy<=SPy+24;
			t<=(others=>'0');
		elsif (estado=S1b) then
			TEx<=VEx-8;
			TEy<=VEy+24;
			t<=(others=>'0');
		elsif (estado=S2a) then
			TEx<=(SPx+24)+(velocidadX*t);
			TEy<="00"&(SPy+24-velocidadY*t+t*t(7 downto 0));
			t<=t+1;
		elsif (estado=S2b) then
			TEx<=(VEx-9)-(velocidadX*t);
			TEy<="00"&(VEy+24-velocidadY*t+t*t(7 downto 0));			
			t<=t+1;
		else
			t<=(others=>'0');
		end if;
	end if;
end process;

-->>> Proceso de obtenci�n de bits en serie en data
process(clkTecl)
begin
	if (clkTecl'event and clkTecl='0') then
		data<=data(9 downto 0) & bitSerie;
	end if;
end process;

-->>> Proceso que valida un valor del teclado
process(reset,clkTecl,contador,estado)
begin
	if (reset='1') then
		tecladoValido<='0';
		dataOk<="00000000";
		dataAnt<="00000000";
		contador<="0000"; -- indica el ciclo por el que vamos. Seg�n el ciclo el valor bitSerie significar� una cosa u otra.
								-- en este caso bitSerie en C1=start, en C2-C9=dato, en C10,C11=paridad,stop
	elsif (clkTecl'event and clkTecl='0') then
		if (estado=S1a or estado=S1b) then
			if (contador="1010") then -- si estamos en C10 tenemos ya el dato en data, porque han pasado los ciclos C2-C9
				dataOk<=data(9 downto 2); -- ...preparamos dataOk para poder mostrar la tecla pulsada por el 7seg en el C11
				dataAnt<=data(9 downto 2); -- ...preparamos dataAnt para poder mostrar la tecla pulsada por el 7seg en los ciclos C1-C10
				contador<="0000";  -- pasamos a C11
				tecladoValido<='1';
			else -- si no estamos en C10...
				dataOk<=dataAnt; -- ...preparamos dataOk para poder mostrar la tecla pulsada por el 7seg en los ciclos siguientes (C2-C11)
				contador<=contador+1; -- ...aumentamos contador
				tecladoValido<='0';
			end if;
		else 
			dataOk<=(others=>'0');
		end if;
	end if;
end process;
			
end vgacore_arch;
